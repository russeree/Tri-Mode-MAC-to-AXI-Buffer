/* Define Simulation */
`define _SIMULATION
/* Verbose debugging */
// `define _dbg_verbose 1
/* Define RST_HOLD and DELAY values relative to timescale */ 
`define _RST_DLY #50
`define _RST_HLD #100
/* BOOLEAN TYPES */ 
`define _true  1'b1
`define _false 1'b0 