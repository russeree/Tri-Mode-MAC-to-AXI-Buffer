/* Define Simulation */
`define _SIMULATION
/* Define RST_HOLD and DELAY values relative to timescale */ 
`define _RST_DLY #50
`define _RST_HLD #100
/* BOOLEAN TYPES */ 
`define _true  1'b1
`define _false 1'b0 